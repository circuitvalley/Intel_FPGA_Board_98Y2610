`timescale 1ns/1ns

module pin_uart_top_tb;
		
pin_uart_top pin_uart_top_ins();
endmodule